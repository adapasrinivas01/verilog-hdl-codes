// port and module
module adder(input a,b,output sum,carry); 
  // or input a,b;
  //    output sum,carrry;
endmodule

// port is the declaration of input and output for the module (a,b,sum,carry)
// module is the basic building block of verilog and it performs specific function
  
